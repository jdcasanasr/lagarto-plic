`define ID_NO_INTERRUPT             32'd0
`define PRIORITY_NEVER_INTERRUPT    32'b0

// ToDo: Define remaining ID's.
`define ID_PLIC                     32'd1
`define ID_JTAG                     32'd2
`define ID_GPIO0                    32'd3
`define ID_GPIO1                    32'd4
`define ID_GPIO2                    32'd5
`define ID_SPI0                     32'd6
`define ID_SPI1                     32'd7
`define ID_DDR                      32'd8
`define ID_DMA                      32'd9
`define ID_UART0                    32'd10
`define ID_UART1                    32'd11
`define ID_UART2                    32'd12
`define TIMER0                      32'd13
`define TIMER1                      32'd14
`define TIMER2                      32'd15

// ToDo: Define proper priorities.
`define PRIORITY_PLIC               32'd1
`define PRIORITY_JTAG               32'd2
`define PRIORITY_GPIO0              32'd3
`define PRIORITY_GPIO1              32'd4
`define PRIORITY_GPIO2              32'd5
`define PRIORITY_SPI0               32'd6
`define PRIORITY_SPI1               32'd7
`define PRIORITY_DDR                32'd8
`define PRIORITY_DMA                32'd9
`define PRIORITY_UART0              32'd10
`define PRIORITY_UART1              32'd11
`define PRIORITY_UART2              32'd12
`define PRIORITY_TIMER0             32'd13
`define PRIORITY_TIMER1             32'd14
`define PRIORITY_TIMER2             32'd15